Stadt
knight
953
266
100
100
10
120
2
100
100
0
100
1
100
100
0
100
1
5
1
1
1
1
1
1
1
1
1
