Haus
archer
950
400
100
100
0
100
1
100
100
0
100
1
100
100
0
100
1
0
1
1
1
1
1
1
1
1
1
